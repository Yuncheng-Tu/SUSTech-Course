module ARM(
    input CLK,
    input Reset,
    input [31:0] Instr,
    input [31:0] ReadData,

    output MemWrite,
    output [31:0] PC,
    output [31:0] ALUResult,
    output [31:0] WriteData
); 
    wire PCSrc;
    wire [31:0] Result, PC, PC_Plus_4;
    wire Busy;
    
    ProgramCounter u_ProgramCounter(
    	.CLK       (CLK       ),
        .Reset     (Reset     ),
        .PCSrc     (PCSrc     ),
        .Result    (Result    ),
        .Busy(Busy),
        .PC        (PC        ),
        .PC_Plus_4 (PC_Plus_4 )
    );


    wire [3:0] ALUFlags;
    
    wire MemtoReg;
    wire MemWrite;
    wire ALUSrc;
    wire [1:0] ImmSrc;
    wire RegWrite;

    wire [2:0] RegSrc;
    wire [1:0] ALUControl;
    //MCycle
    wire M_Start;
    wire MCycleOp;
    wire Mwrite;
    wire [31:0] M_result;
    
    wire done;//���ڶ����ڳ˳��������ˣ�Mwrite����д��
    ControlUnit u_ControlUnit(
    	.Instr      (Instr      ),
        .ALUFlags   (ALUFlags   ),
        .CLK        (CLK        ),
      //  .done(done),
        .MemtoReg   (MemtoReg   ),
        .MemWrite   (MemWrite   ),
        .ALUSrc     (ALUSrc     ),
        .ImmSrc     (ImmSrc     ),
        .RegWrite   (RegWrite   ),
        .RegSrc     (RegSrc     ),
        .ALUControl (ALUControl ),
        .PCSrc      (PCSrc      ),
        .M_Start(M_Start),
        .MCycleOp(MCycleOp),
        .Mwrite(Mwrite)
    );
    

    wire [31:0] Src_A, Src_B, RD2,RD1;
//R F
    wire [3:0] RA1;   assign RA1 = (RegSrc[2])?(Instr[11:8]):((RegSrc[0])?(4'd15):(Instr[19:16]));
    wire [3:0] RA2;   assign RA2 = (RegSrc[2])?(Instr[3:0]):((RegSrc[1])?(Instr[15:12]):(Instr[3:0]));
    wire [3:0] RA3;   assign RA3 = (RegSrc[2])?(Instr[19:16]):(Instr[15:12]);
    
    wire [31:0] PC_Plus_8;
    assign PC_Plus_8 = PC_Plus_4 + 32'd4;
    RegisterFile u_RegisterFile(
    	.CLK (CLK ),
        .WE3 (RegWrite & (~Busy) ),//����һ��~busy, only write when finish multicycle
        .A1  (RA1  ),
        .A2  (RA2  ),
        .A3  (RA3  ),
        .WD3 (Result ),
        .R15 ( PC_Plus_8),
        .RD1 (RD1),
        .RD2 (RD2 )
    );
    
    assign WriteData = RD2;
// Shifter and Extend
    wire [31:0] ExtImm;
    wire [31:0] shift_output;
    assign Src_B = (ALUSrc) ? (ExtImm ): (shift_output);//�Ƿ���λ�Ĵ���������չ������
    assign Src_A= RD1;
    Shifter u_Shifter(
    	.Sh     (Instr[6:5] ),
        .Shamt5 (Instr[11:7] ),
        .ShIn   (RD2   ),
        .ShOut  (shift_output )
    );
    
    Extend u_Extend(
    	.ImmSrc   (ImmSrc   ),
        .InstrImm (Instr[23:0] ),
        .ExtImm   (ExtImm   )
    );
 ////   
    ALU u_ALU(
    	.Src_A      (Src_A      ),
        .Src_B      (Src_B      ),
        .ALUControl (ALUControl ),
        .ALUResult  (ALUResult  ),
        .ALUFlags   (ALUFlags   )
    );
    // RESULT To WD3
    assign Result = (RegSrc[2])?(M_result):((MemtoReg)?(ReadData):(ALUResult));//Mwrite��RegSrc[2]�ǲ���һ���ģ���
        MCycle     #(.width(32))    u_MCycle(
         .CLK(CLK),   // Connect to CPU clock
         .RESET(Reset), // Connect to the reset of the ARM processor.
         .Start(M_Start), // Multi-cycle Enable. The control unit should assert this when MUL or DIV instruction is detected.
         .MCycleOp(MCycleOp), // Multi-cycle Operation. "0" for unsigned multiplication, "1" for unsigned division. Generated by Control unit.
         .Operand1(RD1), // Multiplicand / Dividend
         .Operand2(RD2), // Multiplier / Divisor
         .Result(M_result),  //For MUL, assign the lower-32bits result; For DIV, assign the quotient.
         .Busy(Busy)
    );
endmodule